/*
plyr.v :: player file
*/

module othello

pub fn plyr_henlo() {
	println('aoeu from plyr.v')
}
