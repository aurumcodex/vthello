/*
util.v :: utility file
*/

module othello

pub fn henlo() {
	println('henlo from util.v file')
}
