/*
game.v :: main game logic file
*/

module othello

pub fn game() {
	println('game logic ¯\\_(ツ)_/¯')
}
