/*
algo.v :: algorithm file
*/

module othello

pub fn algo() {
	println('the algo file is where the alpha_beta / negamax / rng move functions would go')
}
