/*
eval.v :: evaluation file
*/

module othello

pub fn eval() {
	println('eval shenanigans')
}
