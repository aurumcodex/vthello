/*
bot.v  :: bot file
*/

module othello

pub fn bot() {
	println('bot logic stuff')
}
