/*
move.v :: moves file
*/

module othello

pub fn move() {
	println('move file says hai')
}
